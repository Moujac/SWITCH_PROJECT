library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use ieee.std_logic_unsigned.all;
use work.switch_pkg.all;

entity mac_controller is
    port(
        clk : in std_logic;
        reset : in std_logic;

        -- Input signals should be active until ack/out is received

        -- Port 0
        macc_in_p0 : in mac_input;
        macc_out_p0 : out mac_output;
        
        -- Port 1
        macc_in_p1 : in mac_input;
        macc_out_p1 : out mac_output;

        -- Port 2
        macc_in_p2 : in mac_input;
        macc_out_p2 : out mac_output;

         -- Port 3
         macc_in_p3 : in mac_input;
        macc_out_p3 : out mac_output;
    );
end mac_controller;

architecture mac_controller_arch of mac_controller is

    -- Make sure multiple requests dont get throught when only one is made in reality
    -- Need to cleate a timeout for mac table

    -- BRAM for MAC table, 8k entries, should be able to read/write in a single cycle by use of duel port
    -- 000 = no port, 001 = port 0 ...
    type mem is array (8191 downto 0) of std_logic_vector(42 downto 0);
    signal mac_table : mem := (others => (others => '0'));
    signal addr_dst, addr_dst_next, addr_src, addr_src_next : std_logic_vector(12 downto 0) := (others => '0');

    -- State machine, who has mem access
    type state_type1 is (P0, P1, P2, P3, NONE);
    signal state_access, state_access_next : state_type1 := NONE;

    -- State machine, who has priority
    type state_type2 is (P0, P1, P2, P3);
    signal state_rr, state_rr_next : state_type2 := P0;

    -- Temp value for hashing, depends on who has access
    signal mac_dst_temp, mac_src_temp : std_logic_vector(47 downto 0);
    signal mac_dst_temp16, mac_src_temp16 : std_logic_vector(15 downto 0);

    -- Counters for timeout
    signal addr_count : std_logic_vector(12 downto 0) := (others => '0');
     -- Should be enough for 100 MHz clock, around 3 hr for overflow, logic for overflow? 
    signal time_count : std_logic_vector(39 downto 0) := (others => '0');

begin
    -- Combinational logic
    -- Can maybe rework so more logic is in combinational part
    process(all) -- VHDL 2008 or above
    begin
        -- Keep val if no change
        state_rr_next <= state_rr;
        state_access_next <= state_access;
        addr_dst_next <= addr_dst;
        addr_src_next <= addr_src;
        -- Maybe redundant
        mac_dst_temp <= (others => '0');
        mac_src_temp <= (others => '0');
        -- Handle who has access, RR based
        -- Prio only changes if highest prio gets its turn!!!
        case state_rr is
            when P0 =>
                if macc_in_p0.req = '1' then
                    state_rr_next <= P1;
                    state_access_next <= P0;
                    mac_dst_temp <= macc_in_p0.mac_dst;
                    mac_src_temp <= macc_in_p0.mac_src;
                elsif macc_in_p1.req = '1' then
                    state_access_next <= P1;
                    mac_dst_temp <= macc_in_p1.mac_dst;
                    mac_src_temp <= macc_in_p1.mac_src;
                elsif macc_in_p2.req = '1' then
                    state_access_next <= P2;
                    mac_dst_temp <= macc_in_p2.mac_dst;
                    mac_src_temp <= macc_in_p2.mac_src;
                elsif macc_in_p3.req = '1' then
                    state_access_next <= P3;
                    mac_dst_temp <= macc_in_p3.mac_dst;
                    mac_src_temp <= macc_in_p3.mac_src;
                else 
                    state_access_next <= NONE;
                end if;
            when P1 =>
                if macc_in_p1.req = '1' then
                    state_rr_next <= P2;
                    state_access_next <= P1;
                    mac_dst_temp <= macc_in_p1.mac_dst;
                    mac_src_temp <= macc_in_p1.mac_src;
                elsif macc_in_p2.req = '1' then
                    state_access_next <= P2;
                    mac_dst_temp <= macc_in_p2.mac_dst;
                    mac_src_temp <= macc_in_p2.mac_src;
                elsif macc_in_p3.req = '1' then
                    state_access_next <= P3;
                    mac_dst_temp <= macc_in_p3.mac_dst;
                    mac_src_temp <= macc_in_p3.mac_src;
                elsif macc_in_p0.req = '1' then
                    state_access_next <= P0;
                    mac_dst_temp <= macc_in_p0.mac_dst;
                    mac_src_temp <= macc_in_p0.mac_src;
                else 
                    state_access_next <= NONE;
                end if;
            when P2 =>
                if macc_in_p2.req = '1' then
                    state_rr_next <= P3;
                    state_access_next <= P2;
                    mac_dst_temp <= macc_in_p2.mac_dst;
                    mac_src_temp <= macc_in_p2.mac_src;
                elsif macc_in_p3.req = '1' then
                    state_access_next <= P3;
                    mac_dst_temp <= macc_in_p3.mac_dst;
                    mac_src_temp <= macc_in_p3.mac_src;
                elsif macc_in_p0.req = '1' then
                    state_access_next <= P0;
                    mac_dst_temp <= macc_in_p0.mac_dst;
                    mac_src_temp <= macc_in_p0.mac_src;
                elsif macc_in_p1.req = '1' then
                    state_access_next <= P1;
                    mac_dst_temp <= macc_in_p1.mac_dst;
                    mac_src_temp <= macc_in_p1.mac_src;
                else 
                    state_access_next <= NONE;
                end if;
            when P3 =>
                if macc_in_p3.req = '1' then
                    state_rr_next <= P0;
                    state_access_next <= P3;
                    mac_dst_temp <= macc_in_p3.mac_dst;
                    mac_src_temp <= macc_in_p3.mac_src;
                elsif macc_in_p0.req = '1' then
                    state_access_next <= P0;
                    mac_dst_temp <= macc_in_p0.mac_dst;
                    mac_src_temp <= macc_in_p0.mac_src;
                elsif macc_in_p1.req = '1' then
                    state_access_next <= P1;
                    mac_dst_temp <= macc_in_p1.mac_dst;
                    mac_src_temp <= macc_in_p1.mac_src;
                elsif macc_in_p2.req = '1' then
                    state_access_next <= P2;
                    mac_dst_temp <= macc_in_p2.mac_dst;
                    mac_src_temp <= macc_in_p2.mac_src;
                else 
                    state_access_next <= NONE;
                end if;
        end case;
        -- Handle hashing, depends on who has access
        -- Simple XOR hashing, maybe not good enough spread
        mac_dst_temp16 <=   mac_dst_temp(47 downto 32) xor mac_dst_temp(31 downto 16) xor 
                            mac_dst_temp(15 downto 0);
        addr_dst_next <=    mac_dst_temp16(12 downto 0);
        mac_src_temp16 <=   mac_src_temp(47 downto 32) xor mac_src_temp(31 downto 16) xor 
                            mac_src_temp(15 downto 0);
        addr_src_next <=    mac_src_temp16(12 downto 0);
    end process;

    -- Sequential logic
    process(clk, reset)
    begin
        if reset = '1' then
            state_access <= NONE;
            state_rr <= P0;
            addr_dst <= (others => '0');
            addr_src <= (others => '0');
            addr_count <= (others => '0');
            time_count <= (others => '0');
        elsif rising_edge(clk) then
            --  Reg update
            state_access <= state_access_next;
            state_rr <= state_rr_next;
            addr_dst <= addr_dst_next;
            addr_src <= addr_src_next;
            time_count <= time_count + 1;
            -- Default output vals
            ack_p0 <= '0';
            ack_p1 <= '0';
            ack_p2 <= '0';
            ack_p3 <= '0';
            out_p0 <= (others => '0');
            out_p1 <= (others => '0');
            out_p2 <= (others => '0');
            out_p3 <= (others => '0');
            -- Handle mem access logic
            case state_access is
                when P0 =>
                    macc_in_p0.outt <= mac_table(to_integer(unsigned(addr_dst)));
                    macc_in_p0.ack <= '1';
                    mac_table(to_integer(unsigned(addr_src))) <= "001" & time_count;
                when P1 =>
                    macc_in_p1.outt <= mac_table(to_integer(unsigned(addr_dst)));
                    macc_in_p1.ack <= '1';
                    mac_table(to_integer(unsigned(addr_src))) <= "010" & time_count;
                when P2 =>
                    macc_in_p2.outt <= mac_table(to_integer(unsigned(addr_dst)));
                    macc_in_p2.ack <= '1';
                    mac_table(to_integer(unsigned(addr_src))) <= "011" & time_count;
                when P3 =>
                    macc_in_p3.outt <= mac_table(to_integer(unsigned(addr_dst)));
                    macc_in_p3.ack <= '1';
                    mac_table(to_integer(unsigned(addr_src))) <= "100" & time_count;
                when NONE =>
                    -- Delete old entries, while memory access is idle
                    addr_count <= addr_count + 1;
                    -- Check if entry is older than 5 minutes at 100 MHz
                    -- 5 minutes = 3000000000 cycles
                    if time_count - mac_table(to_integer(unsigned(addr_count)))(39 downto 0) > x"B2D0000000" then
                        mac_table(to_integer(unsigned(addr_count))) <= (others => '0');
                    end if;
            end case;
        end if;
    end process;
end architecture; 